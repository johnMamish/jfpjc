/**
 * Jpeg requires us to stuff bytes following ff with a 00.
 *
 * This module does that; it needs to handle 32-bit writes, which decreases its efficiency quite a bit.
 */

module bytestuffer();


endmodule
